module Initializer(
    input
    output
);

always_comb begin

end

always_ff @(posedge i_clk or negedge i_rst_n) begin

end

endmodule