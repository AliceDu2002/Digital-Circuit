module RsaPrep(
    input [255:0] N;
    input [255:0] a;
    input [255:0] b;
    input input_ready;
    input [7:0] k;
    output [255:0] m;
    output output_ready;
);

endmodule